module silly (input  logic a, b, c, output logic y);
   
   
   
endmodule
